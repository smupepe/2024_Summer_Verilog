`timescale 1ns/10ps
`define T_CLK 10

module tb_half_adder();
reg din_a;
reg din_b;
wire sum;
wire c_out;

half_adder u_half_adder(
    .din_a(din_a),
    .din_b(din_b),
    .sum(sum),
    .c_out(c_out)
);

initial begin
    din_a = 1'b0;
    din_b = 1'b0;

    #(`T_CLK*1) din_b = 1'b1;
    #(`T_CLK*1) din_a = 1'b1;
               din_b = 1'b0;
    #(`T_CLK*1) din_b = 1'b1;
    #(`T_CLK*1) $stop;
end

endmodule